
Library IEEE;
use IEEE.std_logic_1164.ALL;

Architecture packet_divider_arch of packet_divider is
	begin
		-- create a funtion that divide the packet into symbols
	end architecture;