library IEEE;
use ieee.srd_logic_1164.all;

Entity encoder_ent is
	port( s_id1, s_id2 : in )