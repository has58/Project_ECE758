library IEEE;
use IEEE.std_logic_1164.ALL;


Package network_coding is
	function pack_sym( signal P1, P2 :  in std_logic_vector (63 downto );)
			returen 
