ENtity trial is
	port (a : in symbol;
		b : in packet);
end entity;