-- Author: Haider Ali Siddiquee
-- date : 4/19/2019
-- time 3:21:15 AM
-- package_net_body.vhd
-- contain all the function/proceture definations inside the package

