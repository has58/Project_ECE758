Library IEEE;
use IEEE.std_logic_1164.ALL;

-- Here pac1 and pac2 are two packets
--sym_id1 and sym_id2 are two symbol with their IDs 
-- con_sig is a control signal that control the incoming packet toward the packet divider
Entity packet_divider_ent is 
	port( Pac1, Pac2 : in std_logic_vector (63 downto 0);
		sym_id2, sym_id1 : out std_logic_vector (11 downto 0);
		con_sig : out bit;
		clk : in bit );
end entity; 
